-- heavy citation to Kent Jones's MIPS datapath
library IEEE;
use IEEE.STD_LOGIC_1164.all; 
use IEEE.NUMERIC_STD.all;
use IEEE.math_real.all;
use work.fixed_float_types.all;
use work.float_pkg.all;
use work.fixed_pkg.all;
use IEEE.STD_LOGIC_UNSIGNED.all;

entity control_unit is 
port(instr: in std_logic_vector(63 downto 0) := (others=> '0');
     readBit, writeBit: out std_logic;
     instr_type: out std_logic_vector(1 downto 0) := (others=> '0');
     alucontrol: out std_logic_vector(4 downto 0):= (others=> '0'));
end;

architecture behave of control_unit is
begin 
    instr_type <= instr(63 downto 62);
    alucontrol <= instr(61 downto 57);

    --Set readbit
    with instr(61 downto 57) select readBit <=
        '1' when "01000",
        '0' when others;
    
    --Set writeBit
    with instr(61 downto 57) select writeBit <=
        '1' when "01001",
        '0' when others;
end;
